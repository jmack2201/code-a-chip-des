`timescale 1ns/1ps
module init_perm (
    input [63:0] init_p_box_i,
    output [63:0] init_p_box_o 
);
    assign init_p_box_o[63] = init_p_box_i[57];
    assign init_p_box_o[62] = init_p_box_i[49];
    assign init_p_box_o[61] = init_p_box_i[41];
    assign init_p_box_o[60] = init_p_box_i[33];
    assign init_p_box_o[59] = init_p_box_i[25];
    assign init_p_box_o[58] = init_p_box_i[17];
    assign init_p_box_o[57] = init_p_box_i[9];
    assign init_p_box_o[56] = init_p_box_i[1];
    assign init_p_box_o[55] = init_p_box_i[59];
    assign init_p_box_o[54] = init_p_box_i[51];
    assign init_p_box_o[53] = init_p_box_i[43];
    assign init_p_box_o[52] = init_p_box_i[35];
    assign init_p_box_o[51] = init_p_box_i[27];
    assign init_p_box_o[50] = init_p_box_i[19];
    assign init_p_box_o[49] = init_p_box_i[11];
    assign init_p_box_o[48] = init_p_box_i[3];
    assign init_p_box_o[47] = init_p_box_i[61];
    assign init_p_box_o[46] = init_p_box_i[53];
    assign init_p_box_o[45] = init_p_box_i[45];
    assign init_p_box_o[44] = init_p_box_i[37];
    assign init_p_box_o[43] = init_p_box_i[29];
    assign init_p_box_o[42] = init_p_box_i[21];
    assign init_p_box_o[41] = init_p_box_i[13];
    assign init_p_box_o[40] = init_p_box_i[5];
    assign init_p_box_o[39] = init_p_box_i[63];
    assign init_p_box_o[38] = init_p_box_i[55];
    assign init_p_box_o[37] = init_p_box_i[47];
    assign init_p_box_o[36] = init_p_box_i[39];
    assign init_p_box_o[35] = init_p_box_i[31];
    assign init_p_box_o[34] = init_p_box_i[23];
    assign init_p_box_o[33] = init_p_box_i[15];
    assign init_p_box_o[32] = init_p_box_i[7];
    assign init_p_box_o[31] = init_p_box_i[56];
    assign init_p_box_o[30] = init_p_box_i[48];
    assign init_p_box_o[29] = init_p_box_i[40];
    assign init_p_box_o[28] = init_p_box_i[32];
    assign init_p_box_o[27] = init_p_box_i[24];
    assign init_p_box_o[26] = init_p_box_i[16];
    assign init_p_box_o[25] = init_p_box_i[8];
    assign init_p_box_o[24] = init_p_box_i[0];
    assign init_p_box_o[23] = init_p_box_i[58];
    assign init_p_box_o[22] = init_p_box_i[50];
    assign init_p_box_o[21] = init_p_box_i[42];
    assign init_p_box_o[20] = init_p_box_i[34];
    assign init_p_box_o[19] = init_p_box_i[26];
    assign init_p_box_o[18] = init_p_box_i[18];
    assign init_p_box_o[17] = init_p_box_i[10];
    assign init_p_box_o[16] = init_p_box_i[2];
    assign init_p_box_o[15] = init_p_box_i[60];
    assign init_p_box_o[14] = init_p_box_i[52];
    assign init_p_box_o[13] = init_p_box_i[44];
    assign init_p_box_o[12] = init_p_box_i[36];
    assign init_p_box_o[11] = init_p_box_i[28];
    assign init_p_box_o[10] = init_p_box_i[20];
    assign init_p_box_o[9] = init_p_box_i[12];
    assign init_p_box_o[8] = init_p_box_i[4];
    assign init_p_box_o[7] = init_p_box_i[62];
    assign init_p_box_o[6] = init_p_box_i[54];
    assign init_p_box_o[5] = init_p_box_i[46];
    assign init_p_box_o[4] = init_p_box_i[38];
    assign init_p_box_o[3] = init_p_box_i[30];
    assign init_p_box_o[2] = init_p_box_i[22];
    assign init_p_box_o[1] = init_p_box_i[14];
    assign init_p_box_o[0] = init_p_box_i[6];
endmodule