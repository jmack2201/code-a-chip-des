module final_perm (
    input [1:64] final_p_box_i,
    output [1:64] final_p_box_o 
);
    assign final_p_box_o[1] = final_p_box_i[40];
    assign final_p_box_o[2] = final_p_box_i[8];
    assign final_p_box_o[3] = final_p_box_i[48];
    assign final_p_box_o[4] = final_p_box_i[16];
    assign final_p_box_o[5] = final_p_box_i[56];
    assign final_p_box_o[6] = final_p_box_i[24];
    assign final_p_box_o[7] = final_p_box_i[64];
    assign final_p_box_o[8] = final_p_box_i[32];
    assign final_p_box_o[9] = final_p_box_i[39];
    assign final_p_box_o[10] = final_p_box_i[7];
    assign final_p_box_o[11] = final_p_box_i[47];
    assign final_p_box_o[12] = final_p_box_i[15];
    assign final_p_box_o[13] = final_p_box_i[55];
    assign final_p_box_o[14] = final_p_box_i[23];
    assign final_p_box_o[15] = final_p_box_i[63];
    assign final_p_box_o[16] = final_p_box_i[31];
    assign final_p_box_o[17] = final_p_box_i[38];
    assign final_p_box_o[18] = final_p_box_i[6];
    assign final_p_box_o[19] = final_p_box_i[46];
    assign final_p_box_o[20] = final_p_box_i[14];
    assign final_p_box_o[21] = final_p_box_i[54];
    assign final_p_box_o[22] = final_p_box_i[22];
    assign final_p_box_o[23] = final_p_box_i[62];
    assign final_p_box_o[24] = final_p_box_i[30];
    assign final_p_box_o[25] = final_p_box_i[37];
    assign final_p_box_o[26] = final_p_box_i[5];
    assign final_p_box_o[27] = final_p_box_i[45];
    assign final_p_box_o[28] = final_p_box_i[13];
    assign final_p_box_o[29] = final_p_box_i[53];
    assign final_p_box_o[30] = final_p_box_i[21];
    assign final_p_box_o[31] = final_p_box_i[61];
    assign final_p_box_o[32] = final_p_box_i[29];
    assign final_p_box_o[33] = final_p_box_i[36];
    assign final_p_box_o[34] = final_p_box_i[4];
    assign final_p_box_o[35] = final_p_box_i[44];
    assign final_p_box_o[36] = final_p_box_i[12];
    assign final_p_box_o[37] = final_p_box_i[52];
    assign final_p_box_o[38] = final_p_box_i[20];
    assign final_p_box_o[39] = final_p_box_i[60];
    assign final_p_box_o[40] = final_p_box_i[28];
    assign final_p_box_o[41] = final_p_box_i[35];
    assign final_p_box_o[42] = final_p_box_i[3];
    assign final_p_box_o[43] = final_p_box_i[43];
    assign final_p_box_o[44] = final_p_box_i[11];
    assign final_p_box_o[45] = final_p_box_i[51];
    assign final_p_box_o[46] = final_p_box_i[19];
    assign final_p_box_o[47] = final_p_box_i[59];
    assign final_p_box_o[48] = final_p_box_i[27];
    assign final_p_box_o[49] = final_p_box_i[34];
    assign final_p_box_o[50] = final_p_box_i[2];
    assign final_p_box_o[51] = final_p_box_i[42];
    assign final_p_box_o[52] = final_p_box_i[10];
    assign final_p_box_o[53] = final_p_box_i[50];
    assign final_p_box_o[54] = final_p_box_i[18];
    assign final_p_box_o[55] = final_p_box_i[58];
    assign final_p_box_o[56] = final_p_box_i[26];
    assign final_p_box_o[57] = final_p_box_i[33];
    assign final_p_box_o[58] = final_p_box_i[1];
    assign final_p_box_o[59] = final_p_box_i[41];
    assign final_p_box_o[60] = final_p_box_i[9];
    assign final_p_box_o[61] = final_p_box_i[49];
    assign final_p_box_o[62] = final_p_box_i[17];
    assign final_p_box_o[63] = final_p_box_i[57];
    assign final_p_box_o[64] = final_p_box_i[25];

endmodule
